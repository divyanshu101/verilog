module frst();

$display("hellow");
endmodule
